1.7.14 - Resonant Circuits, Figure 1.106
* 
* Author : Nicolas Misbert 
* Source : Art Of Electronics, Third Edition
*   Paul Horowitz
*   Winfield Hill
*
vin in 0 pulse(0.0V 2.0V 2ms) ac 1.0 dc 0.0
r1 in out 10k
c1 out 0 0.1u
l1 out 0 0.2k

.control 
tran 0.1ms 10ms 0.0ms 0.2ms
ac dec 10 1.0Hz 10kHz
plot (v(out)/v(in)) xlog
.endc
.end