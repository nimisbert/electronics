* Circuit :
* Ideal Colpitts Oscillator
Ec C 0 table {2.5*V(E)} (0.5 0.5 14.5 14.5) ; Low (0.5V) High (14.5V) limits
R1 C S 47
C1 S E 30p
C2 E 0 30p
Rl E 0 1Meg
L1 S 0 220n
.ic V(E) = 2V
.tran .1ns 150ns 0n .1ns
.probe
.end