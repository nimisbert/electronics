* Circuit :
* Exemple avec OP
V1 1 0 DC=1
V2 2 0 DC=2
R1 1 3 3.3k
R2 2 3 6.8k
R3 3 0 4.7k
.op
.end
* +----R1----+
* |          |
* |   +--R2--+---+
* |   |      |   |
* V1  V2     R3  S
* |   |      |   |
* +---+-gnd--+---+