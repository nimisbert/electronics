2.2.4 - Emitter followers as voltage regulators, Figure 2.20.
* 
* Author : Nicolas Misbert 
* Source : Art Of Electronics, Third Edition
*   Paul Horowitz
*   Winfield Hill
*
.model ZEN D (BV=10 IBV=17m) 

vin in 0 sin(22.5 2.5 20) dc 0.0
r1 in out 1k
d1 0 out ZEN

.control 
delete all
tran 200us 200ms 0ms 1ms
plot v(in) v(out)
.endc
.end