4.1.2 - Pulse-Generator III, Figure 2.13.A.
* 
* Author : Nicolas Misbert 
* Source : Art Of Electronics, Third Edition
*   Paul Horowitz
*   Winfield Hill
*
.model QMOD NPN (level=4 IS=1.6e-16)

vsupply 1  0 dc 5V
vlogic  in 0
r7      1  2 1k 
r6      in 3 25k
q4      2 3 4 QMOD IC=0.6
r9      4 0 20
r8      1 out 1k
q5      out 2 4 QMOD IC=0.6

.control 
dc vlogic 0.0 3.3 +0.1
plot v(in) v(out)
.endc
.end