1.6.7 - Inductive loads and diode protection, Figure 1.83.
* 
* Author : Nicolas Misbert 
* Source : Art Of Electronics, Third Edition
*   Paul Horowitz
*   Winfield Hill
*
.model SWITCH sw( VT=1.0 VH=0.0 )
.model ROLLBACK D( IS=18.8n BV=0.1 IBV=5.00u )

vs supply  0 dc 1.0
vl control 0 dc 0.0 pulse(0.0V 1.0V 2ms)
l1 supply  1 100n
s1 1 0 control 0 SWITCH

l2 supply  2 100n 
d2 2 supply ROLLBACK
s2 2 0 control 0 SWITCH

l3 supply 3 100n
r3 supply 4 100
c3 4 3 0.05u
s3 3 0 control 0 SWITCH

.control
delete all
tran 0.1ms 2.101ms 2.0999ms 0.00001ms
let kick = v(1)
let rollback = v(2)
let snubber = v(3)
plot kick snubber rollback
destroy
.endc 
.end 