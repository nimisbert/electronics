* Circuits with Diodes
* Diode model
.model ID D(Ron=1 Roff=1Meg Vfwd=0 Vrev=75)

* --- Half-wave rectifier --- *
* 1-D|-2
*V1 1 0 SINE(0 3.3 50)
*D1 1 2 ID
*R1 2 0 1k
*.tran 0.06

* --- Full-wave rectifier --- *
*   +-D|1-+1+-D|2-+
* 3-+             +-4
*   +-D|3-+2+-D|4-+
*V2 1 2 SINE(0 10 50)
*D1 0 1 ID
*D2 1 4 ID
*D3 0 2 ID
*D4 2 4 ID
* Vdc = sqrt(2) * Vac (rms)
* Ripple Half-bridge = Iload / f*C
* Ripple Full-bridge = Iload / 2*f*C
*C2 4 0 .002 ; power filtering
*R2 4 0 1k
*.tran 0.10

* --- Center Tapped Full-wave rectifier --- *
* Primary
*V3 1 0 SINE(0 10 50)
*Rv 1 2 10 ; prevent over defined circuit
*L1 2 0 10m
* Secondary
*L2 3 0 10u
*L3 0 4 10u
*D1 3 6 ID
*D2 4 7 ID
*R2 6 7 1k
*K1 L1 L2 L3 1.0

* --- Dual Polarity Split Supply --- *
* Primary
*V3 1 0 SINE(0 10 50)
*Rv 1 2 1 ; prevent over defined circuit
*L1 2 0 1u
* Secondary
*L2 4 0 1
*L3 0 6 1
*D1 3 4 ID
*D2 4 5 ID
*D3 3 6 ID
*D4 6 5 ID
*C1 3 0 1u
*C2 5 0 1u
*K1 L1 L2 L3 1.0
*.tran 0.10

* --- Voltage Multipliers --- *
* --- Cockcroft-Walton CW --- *
* Primary
*V3 1 0 SINE(0 10 50)
*Rv 1 2 1 ; prevent over defined circuit
*L1 2 0 1u
* Secondary
*L2 4 3 1
*L3 3 0 1
*K1 L1 L2 L3 1.0
* CW First Stage
*C1 4 5 1u
*C2 6 0 1u
*D1 0 5 ID
*D2 5 6 ID
* CW Second Stage (Voltage Doubler)
*C3 5 7 1u
*C4 6 8 1u
*D3 6 7 ID
*D4 7 8 ID
* CW Third Stage (Voltage Tripler)
*C5 7 9 1u
*C6 8 10 1u
*D5 8 9 ID
*D6 9 10 ID
* CW Fourth Stage (Voltage Quadrupler)
*C7 9 11 1u
*C8 10 12 1u
*D7 10 11 ID
*D8 11 12 ID
*.tran 0.60

* --- Signal Rectifier --- *
*V1 1 0 pulse (0 3 100u 1n 1n 200u 400u)
*C1 1 2 0.1u
*R1 2 0 100
*D1 2 3 ID
*R2 3 0 100
*.tran 1200u

* --- Signal Rectifier with Voltage Drop Compensation --- *
*V1 1 0 pulse (0 0.5 100u 1n 1n 200u 400u)
*V2 4 0 DC=5
*C1 1 2 100p
*R1 2 3 1k
*D1 3 0 ID
*R2 3 4 1k
*D2 2 5 ID
*R3 5 0 1k
*.tran 1200u

* --- Diode Clamp --- *
* Circuit Figure 1.72
* Clamps above 5.6V
*V1 in 0 SINE(0 10 50)
*V2 3 0 dc 5
*R1 in out 1k
*D1 out 3 ID
*.tran 0.20

* Clamps below -5.6V
*V1 in 0 SINE(0 10 50)
*R1 in out 1k
*D1 3 out ID
*Vc 3 0 dc -5.6
*.tran 0.10

* Circuit Exercice 1.22
* Symetrical clamp from -5.6 to 5.6
*V1 in 0 SINE(0 10 50)
*R1 in out 1k
*DclampP out vcp ID
*DclampM vcm out ID
*VclampP vcp 0 dc 5.6
*VclampM vcm 0 dc -5.6
*.tran 0.10

* --- Diode Clamp --- *
* Circuit Figure 1.78
*V1 in 0 SINE(0 10 50)
*R1 in out 1k
*D1 out 0 ID
*D2 0 out ID
*.tran 0.10

* TODO
* --- Non-Linear elements --- *
* Circuit Figure 1.80 logarithmic converter
*I1 io 0 1 <------ FAIRE RAMPE DE 0.0 A 20.0
*D1 io 0 ID
*.tran 0.10

* TODO
* Circuit Figure 1.84 inductive kick-blocker
*V1 in 0 DC=10
*L1 in out 1u
*D1 out in
** SW **


.probe
.end