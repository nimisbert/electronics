2.2.2.B - Variations on a theme, Figure 2.10.A.
* 
* Author : Nicolas Misbert 
* Source : Art Of Electronics, Third Edition
*   Paul Horowitz
*   Winfield Hill
*
.model QMOD PNP (level=4 IC=0.6)

vsupply 1 0 dc 15.0V
vlogic  2 0 pulse(15.0V 0.0V 2ms) dc 0.0
rb      2 3 3.3k
q1      1 3 4 QMOD
rload   4 0 10k

.control
delete all
tran 0.1ms 10ms 0.0ms 0.2ms
plot v(4) v(2)
.endc
.end 