2.2.4 - Emitter Followers as voltage regulators, Figure 2.21.
* 
* Author : Nicolas Misbert 
* Source : Art Of Electronics, Third Edition
*   Paul Horowitz
*   Winfield Hill
*
.model ZEN D (BV=10 IBV=17m) 
.model QMOD NPN (level=4 IS=1.6e-16)

vin in 0 sin(22.5 2.5 20) dc 0.0
rb in 1 10k
rc in 2 1k
d1 0 1 ZEN
q1 2 1 out QMOD IC=0.6

.control 
delete all
tran 200us 200ms 0ms 1ms
plot v(in) v(out)
.endc
.end