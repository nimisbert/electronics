* Circuit :
* ----R---+---+
* |       |   |
* |       C1  |
* Vin  ---+   L
* |    |  C2  |
* |    Rl |   |
* |    |  |   |
* +-gnd+--+---+
Vin C 0 AC 1
R1 C S 47
C1 S E 30p
C2 E 0 30p
L1 S 0 220n
Rl E 0 1Meg
.ac dec 100 1Meg 10G
.probe
.end