2.2.2.A - Switching circuit examples, Figure 2.9
* 
* Author : Nicolas Misbert 
* Source : Art Of Electronics, Third Edition
*   Paul Horowitz
*   Winfield Hill
*
.model LED D (AREA=3.0 IC=0.2)
.model QMOD NPN (level=4 IC=0.6)

vsupply 1 0 dc 3.3V
vlogic  2 0 pulse(0.0V 3.3V 2ms) dc 0.0
d1      3 1 LED 
rc      3 4 330
rb      2 5 10k
q1      4 5 0 QMOD

.control
delete all
tran 0.1ms 10ms 0.0ms 0.2ms
plot v(2) v(3)
.endc
.end 