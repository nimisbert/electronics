Exercise 1.1
* 
* Source : The Art Of Electronics, 3rd Edition
* Author : Paul Horowitz, Winfield Hill
* Solver : nimisbert
* Brief :
* You have a 5k resistor and a 10k resistor. 
* What's their combined resistance :
* (a) in series and (b) in parallel ?
*

r1 1 2 5k
r2 2 0 10k
i1 0 1 1A

r3 3 0 5k
r4 3 0 10k
i2 0 3 1A

.control
op
echo En fixant I=1A, U=R, la mesure de V donne Req
echo a)
print v(1)
echo b) 
print v(3)

.endc
.end
