* LF411 operational amplifier
* "macromodel" subcircuit
*
* connections:
*    1 -  non-inverting input
*    2 -  inverting input
*    3 -  positive power supply
*    4 -  negative power supply
*    5 -  output
*
.subckt LF411/MC  1 2 3 4 5
*
  c1   11 12 2.801E-12
  c2    6  7 8.000E-12
  css  10 99 3.200E-12
  dc    5 53 dx
  de   54  5 dx
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 3.316E6
+ -3E6 3E6 3E6 -3E6
  ga    6  0 11 12 402.1E-6
  gcm   0  6 10 99 12.72E-9
  iss   3 10 dc 280.0E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   4 11 2.487E3
  rd2   4 12 2.487E3
  ro1   8  5 40
  ro2   7 99 60
  rp    3  4 24.00E3
  rss  10 99 714.3E3
  vb    9  0 dc 0
  vc    3 53 dc 1.100
  ve   54  4 dc .3
  vlim  7  8 dc 0
  vlp  91  0 dc 30
  vln   0 92 dc 30
.model dx D(Is=800.0E-18)
.model jx PJF(Is=30.00E-12 Beta=577.5E-6
+ Vto=-1)
.ends
*$


