2.2.2.B - Variations on a theme, Figure 2.10.B.
* 
* Author : Nicolas Misbert 
* Source : Art Of Electronics, Third Edition
*   Paul Horowitz
*   Winfield Hill
*
.model QPNP PNP (level=4 IC=0.6)
.model QNPN NPN (level=4 IC=0.6)

vsupply 1 0 dc 15.0V
vlogic  2 0 pulse(0.0V 3.3V 2ms 0.01ms 0.01ms 2ms 10.0ms) dc 0.0
r3      1 3 1k
r2      3 4 3.3k
r1      2 5 10k
q2      4 5 0 QNPN
q3      1 3 6 QPNP
rload   6 0 10k

.control
delete all
tran 0.1ms 6ms 0.0ms 0.2ms
plot v(2) v(3) v(6)
.endc
.end