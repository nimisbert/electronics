2.2.2.C - Pulse-Generator - I, Figure 2.11
* 
* Author : Nicolas Misbert 
* Source : Art Of Electronics, Third Edition
*   Paul Horowitz
*   Winfield Hill
*
.model QMOD NPN (level=4 IC=0.6)

vsupply 1 0 dc 5V
vlogic  in 0 pulse(0.0V 3.3V 1ms) dc 0.0
r1      in 2 10k
r2      1 3 1k
q1      3 2 0 QMOD
c1      3 4 10n
r3      1 4 10k
r4      1 out 1k
q2      out 4 0 QMOD

.control 
delete all
tran 0.01ms 1.4ms 0.8ms 0.1ms
plot v(in) v(out) v(4)
.endc
.end