2.2.3.C - Emitter drives switch, Figure 2.15.B.
* 
* Author : Nicolas Misbert 
* Source : Art Of Electronics, Third Edition
*   Paul Horowitz
*   Winfield Hill
*

.model LED D (BV=3.6 IBV=0.5 IS=100pA N=1.679)
.model QMOD NPN (level=4)

vin    supply 0 5.00 ac 1 dc 5.0
vlogic in 0 1.00 ac 1 dc 3.3 pulse(0.0V 3.3V 2ms) 
d1     supply 1 LED
r2     1  4 220
r4     2  3 100
q3     4  3 0 QMOD IC=0.6
q2     supply in 2 QMOD IC=0.6
r3     2  0 10k

.control 
delete all
tran 200us 4ms 0ms 1ms
plot v(supply) v(in) v(4)
.endc
.end