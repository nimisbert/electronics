* Circuit
V1 1 0 1
R1 1 2 1
R2 2 3 3.3
R3 3 4 2.2
R4 4 0 8.2
R5 0 2 4.7
R6 2 4 6.8
.OP
.end