0 - Voltage Divider to test setup
*
* Author : Nicolas Misbert 
* Source : 
*
vin 1 0 dc
r1 1 2 1.0k
r2 2 0 1.0k

.control
delete all
* dc <src> <start> <stop> <step>
dc vin 0.0V 5.0V 1.0V
plot v(1) v(2)
op
destroy
.endc
.end