* Circuit :
* Colpitts Final Model
.include 2N2222.mod
* A
Vcc A 0 DC=15
RB2 A B 150k
RB1 B 0 22k
Cde B 0 100n
Q1 C B E 2N2222
RE E 0 1040
L1 A C 220n
* b
C1 C E 30p
C2 E 0 30p

*.op
.ic V(E) = 2V
.tran 10p 1u .3u 10p
.probe
.end