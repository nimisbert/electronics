0 - Voltage Divier
*
* Author : Nicolas Misbert 
* Source : 
*
v1 1 0 sin(1 1 10) dc 0.0
r1 1 2 1.0k
r2 2 0 1.0k

.control
delete all
run
op
tran 0.1ms 0.1s 0.1ms 0.1ms
plot v(1) v(2)
destroy
.endc
.end