0 - Testing Basic diode model

.model LED D (BV=3.5 IBV=0.5 IS=100pA N=1.679)

vin in 0 1.00 ac 1 dc 0.0
d1  in 1 LED
r1  1 0 220


.control 
delete all
dc vin -10.0 10.0 0.1
plot i(vin) vs v(in) 
.endc
.end